`ifndef AXI_LITE_COMMON_SV
`define AXI_LITE_COMMON_SV

parameter int MAX_VALUE = 255;
parameter int WIDTH = 9;
parameter int COLUMNS_REG_ADDR = 0;
parameter int LINES_REG_ADDR = 4;
parameter int START_REG_ADDR = 8;
parameter int READY_REG_ADDR = 12;

`endif // AXI_LITE_COMMON_SV
